module MEM(
    input  clk,
    input  rst,
    input  [63:0] EX_pc_i,
    output [63:0] MEM_pc_o,
);

endmodule