module ex();


endmodule